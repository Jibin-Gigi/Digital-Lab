`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:45:16 04/15/2024 
// Design Name: 
// Module Name:    AND_Gate 
// Project Name: Logic_Gates
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module AND_Gate(
    input a,
    input b,
    output y
    );

and(y,a,b);
endmodule
